package constant_package is

    constant C_TIMER_MAX : positive := 60 * 100;

end constant_package;