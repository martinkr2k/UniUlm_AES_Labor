library ieee;
use ieee.std_logic_1164.all;

entity light is 
  port (
    x1 : in std_logic;
    x2 : in std_logic;
    f  : out std_logic
  );
end light;

architecture DATAFLOW of light is
  begin 

    f <= (x1 AND not(x2)) OR (not(x1) AND x2);

end DATAFLOW;
