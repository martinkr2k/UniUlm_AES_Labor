library ieee;
use ieee.std_logic_1164.all;

entity fourbit_fa is 
  port (
    sw : in std_logic_vector(9 downto 0);
    ledr : out std_logic_vector(9 downto 0)
  );
end fourbit_fa;


architecture DATAFLOW of fourbit_fa is 
  signal s_ctemp : std_logic_vector(4 downto 0);
  begin 

    FA0 : entity work.fa(DATAFLOW) port map(sw(0), sw(4), s_ctemp(0), ledr(0), s_ctemp(1));
    FA1 : entity work.fa(DATAFLOW) port map(sw(1), sw(5), s_ctemp(1), ledr(1), s_ctemp(2));
    FA2 : entity work.fa(DATAFLOW) port map(sw(2), sw(6), s_ctemp(2), ledr(2), s_ctemp(3));
    FA3 : entity work.fa(DATAFLOW) port map(sw(3), sw(7), s_ctemp(3), ledr(3), s_ctemp(4));
	 
	 s_ctemp(0) <= sw(8);
    ledr(4) <= s_ctemp(4);
	 
end DATAFLOW;