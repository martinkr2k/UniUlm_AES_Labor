package constant_package is

    constant C_POLYNOM : positive := 8;
    constant C_MESSAGE : positive := 32;

end constant_package;